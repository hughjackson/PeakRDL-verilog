{%- macro body(node, offset='', index='') %}
// ============================================================
// Register: {{node.get_rel_path(node.parent).upper()}}
{%- for child in node.fields() %}
//    [{{child.bit_range}}] {{'%20s'%child.get_rel_path(node)}}: hw={{'%-5s'%child.get_property('hw').name}} sw={{'%-5s'%child.get_property('sw').name}} reset=0x{{'%x'%(child.get_property('reset') or 0)}}
{%- endfor %}
// ============================================================
logic                  {{signal(node)}}_decode;
logic                  {{signal(node)}}_sw_wr;
logic                  {{signal(node)}}_sw_rd;
logic [DATA_WIDTH-1:0] {{signal(node)}}_q;

assign {{signal(node)}}_decode = (addr == ({{offset}}));
assign {{signal(node)}}_sw_wr = valid && !read && {{signal(node)}}_decode;
assign {{signal(node)}}_sw_rd = valid &&  read && {{signal(node)}}_decode;

assign {{signal(node)}}_strb{{index}} = {{signal(node)}}_sw_wr;

always_comb begin
    {{signal(node)}}_q[{{node.bit_range}}] = '0;
{%- for child in node.fields() %}
    {{signal(node)}}_q[{{child.bit_range}}] = {{signal(child)}}_q{{index}};
{%- endfor %}
end

// masked version of return data
assign {{signal(node)}}_rdata{{index}} = {{signal(node)}}_sw_rd ? {{signal(node)}}_q : 'b0;

{%- for child in node.fields() %}

// Field: {{child.get_rel_path(node)}} 

{%- if not child.implements_storage %}
    {%- if child.is_hw_writable %}
assign {{signal(child)}}_q{{index}} = {{signal(child)}}_wdata;

    {%- else %}
assign {{signal(child)}}_q{{index}} = {{child.get_property('reset')}};

    {%- endif %}
{%- else %}
always_ff @ (posedge clk, negedge resetn)
    if (~resetn) begin
        {{signal(child)}}_q{{index}} <= {{child.get_property('reset', default=0)}};
    end else begin
        {%- if child.is_sw_writable %}
        // Software write
        if ({{signal(node)}}_sw_wr) begin
        {%- if child.get_property('onwrite') == OnWriteType.wclr %}
            {{signal(child)}}_q{{index}} <= 'b0;
        {%- else %}
            {{signal(child)}}_q{{index}} <= (wdata[{{child.bit_range}}] & mask[{{child.bit_range}}]) | ({{signal(child)}}_q{{index}}[{{child.bit_range}}] & ~mask[{{child.bit_range}}]);
        {%- endif %}
        end
        {%- endif -%}

        {%- if child.is_hw_writable %}
        // Hardware Write
        if ({{signal(child)}}_wr{{index}}) begin
            {{signal(child)}}_q{{index}} <= {{signal(child)}}_wdata{{index}};
        end
        {%- endif -%}

        {%- if child.is_up_counter %}
        // Counter increment
        if ({{signal(child)}}_incr{{index}}) begin
            {{signal(child)}}_q{{index}} <= {{signal(child)}}_q{{index}} + {{get_counter_value(child, index, 'incr')}};
        end
        {%- endif %}
        {%- if child.is_down_counter %}
        // Counter decrement
        if ({{signal(child)}}_decr{{index}}) begin
            {{signal(child)}}_q{{index}} <= {{signal(child)}}_q{{index}} - {{get_counter_value(child, index, 'decr')}};
        end
        {%- endif %}
    end

{%- endif %}

{%- endfor -%}
{%- endmacro %}
